// 4-bit counter RTL code
module down_counter    // Module start declaration
 // Parameter declaration, count signal width set to '4'  
 #(parameter WIDTH=4)  
 ( 
    input logic clk,
    input logic clear, 
    output logic[WIDTH-1:0] count
 );

 // Student to add code for down counter logic

 
endmodule: down_counter  // Module end declaration